`include "rom.v"
module rom_tb();
parameter DW=8,
	  AW=4,
	  DEP=16;
reg               wr,rst;       
reg      [DW-1:0] data;
reg      [AW-1:0] addr;
wire     [DW-1:0] data_out;

rom dut(.rst(rst),
	.wr(wr),
	.data(data),
	.addr(addr),
	.data_out(data_out));
initial begin
rst=1'b1;
#10;
rst=1'b0;
wr=1'b0;
addr=4'd8;
#10;
wr=1'b1;
data=8'b0101_0001;
addr=4'd8;
#10;
wr=1'b0;
#10;
#10;

$finish;
end

always@(data_out) begin
 if (data_out[7]==1'b1 && data_out[5]==1'b1) $display("ROM test is PASSESD!!!");
end

endmodule
