module rr_tb();
reg clk,rstn;
reg [3:0] req;
wire [3:0] grant;
wire [3:0] ack;
round_robin dut(.clk(clk),.rstn(rstn),.req(req),.grant(grant),.ack(ack));

initial begin
clk=1'b1;
forever #5 clk=~clk;
end

initial begin
reset();
if($test$plusargs("priority")) begin
 @(negedge clk);
 req=4'b1100;
 n_delay(10);
 @(negedge clk);
 req=4'b1110;
 n_delay(14);
 @(negedge clk);
 req=4'b1111;
 n_delay(18);
 @(negedge clk);
 req=4'b1000;
 n_delay(5);
end
if($test$plusargs("S0")) begin
@(negedge clk);
req=4'b0101;
n_delay(11); // 4 + 4 cycle for 2 ones and 2 cycle for IDLE case 1 cycle for engedge on another req
 req=4'b1001;
 n_delay(11);
 req=4'b0011;
 n_delay(11);
 req=4'b0001;
 n_delay(6);
end

if($test$plusargs("S1")) begin
@(negedge clk);
req=4'b0110;
n_delay(11); // 4 + 4 cycle for 2 ones and 2 cycle for IDLE case 1 cycle for engedge on another req
 req=4'b1010;
 n_delay(11);
 req=4'b0010;
 n_delay(5);
 req=4'b0001;
 n_delay(7);
 req=4'b0010;
 n_delay(6);
end

if($test$plusargs("S2")) begin
@(negedge clk);
req=4'b1100;
n_delay(11); // 4 + 4 cycle for 2 ones and 1 for ack 1 cycle for IDLE case 1 cycle for engedge on another req
 req=4'b0100;
 n_delay(5);
 req=4'b0001;
 n_delay(7);
 req=4'b0100;
 n_delay(5);
 req=4'b0010;
 n_delay(7);
 req=4'b0100;
 n_delay(6);
end

if($test$plusargs("S3")) begin
@(negedge clk);
 req=4'b1000;
 n_delay(4);
 req=4'b0001;
 n_delay(7);
  req=4'b1000;
 n_delay(5);
 req=4'b0010;
 n_delay(7);
 req=4'b1000;
 n_delay(5);
 req=4'b0100;
 n_delay(7);
 req=4'b1000;
 n_delay(6);
end

//repeat(20) @(negedge clk);
$finish;
end

task reset();
	begin
	rstn=1'b0;
	@(negedge clk);
	rstn=1'b1;
end
endtask
task n_delay(input integer n);
begin
 repeat(n) @(negedge clk);
end
endtask
endmodule
