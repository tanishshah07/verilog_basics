`include "main.v"

module top();
reg clk,rst,in;
wire p,c;

main dut(.p(p),.c(c),.clk(clk),.rst(rst),.in(in));

initial forever #5 clk=~clk;

initial begin
rst=1'b0;
clk=0;
@(negedge clk);
reset();

// test case 4(10)
in=1;
@(negedge clk);
in=0;
@(negedge clk);
@(negedge clk);

//test case 1 (111)
reset();
in=1;
@(negedge clk);
in=1;
@(negedge clk);
in=1;
@(negedge clk);
@(negedge clk);
in=1;
@(negedge clk);

// test case 2(01)
reset();
in=0;
@(negedge clk);
in=1;
@(negedge clk);

// test case 3(00)
reset();
in=0;
@(negedge clk);
in=0;
// test case 4(10)
reset();
in=1;
@(negedge clk);
in=0;
@(negedge clk);
// test case 5(110)
reset();
in=1;
@(negedge clk);
in=1;
@(negedge clk);
in=1;
@(negedge clk);
in=0;
//test for default
dut.state=3'd5;
in=1'b1;
@(negedge clk);
dut.state=3'd5;
in=1'b0;
@(negedge clk);
repeat(10) @(negedge clk);
$finish;



end
task reset();
	begin
	 rst=1;
	 @(negedge clk);
	 rst=0;

	end

endtask



endmodule
