module rr(clk,rstn,);




endmodule
